// Top module
