// Testbench code
