// SystemVerilog code for Hamming Encoder
