// RAID 5 Controller logic
